class axi_sequence extends uvm_sequence #(axi_transaction);
endclass