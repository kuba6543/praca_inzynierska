class axi_agent extends uvm_agent;
  	// declaring agent components
    axi_driver    driver;
    axi_sequencer sequencer;
    axi_monitor   monitor;

	// hold parameter if the agent is slave
    bit is_slave;

  	// UVM automation macros for general components
    `uvm_component_utils(axi_agent)

  	// constructor of AXI agent
    function new (string name, uvm_component parent);
        super.new(name, parent);
    endfunction : new

    // build agent, whether is passive or active
    function void build_phase(uvm_phase phase);
        super.build_phase(phase);
        if(get_is_active() == UVM_ACTIVE) begin
            driver = axi_driver::type_id::create("driver", this);
            sequencer = axi_sequencer::type_id::create("sequencer", this);
        end
        monitor = axi_monitor::type_id::create("monitor", this);
        uvm_config_db#(bit)::set(this, "driver", "is_slave", is_slave);
    endfunction : build_phase

  	// connect driver with sequencer if the agent is active
    function void connect_phase(uvm_phase phase);
        if(get_is_active() == UVM_ACTIVE) begin
        driver.seq_item_port.connect(sequencer.seq_item_export);
    end
    driver.is_slave = this.is_slave;
    endfunction : connect_phase

endclass : axi_agent