`include "axi_agent/axi_sequencer.sv"
`include "axi_agent/axi_driver_slave.sv"
`include "axi_agent/axi_driver_master.sv"
`include "axi_agent/axi_monitor.sv"
`include "axi_agent/axi_agent_slave.sv"
`include "axi_agent/axi_agent_master.sv"
`include "axi_sequence.sv"
`include "axi_transaction.sv"
`include "axi_scoreboard.sv"
`include "axi_enviroment.sv"
`include "axi_test.sv"