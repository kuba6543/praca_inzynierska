class axi_transaction extends uvm_sequence_item;
endclass